module XOR_Gate(
    input wire A,   // First input
    input wire B,   // Second input
    output wire Y   // Output
);

    assign Y = A ^ B; // XOR operation

endmodule
