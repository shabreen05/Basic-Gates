module NOT_Gate(
    input wire A,   // Input
    output wire Y   // Output
);

    assign Y = ~A; // NOT operation

endmodule
